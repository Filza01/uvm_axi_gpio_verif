package gpio_pkg;

    import uvm_pkg::*;
   `include "uvm_macros.svh"
  
   `include "env_gpio/gpio_seq_item.sv"
   `include "env_gpio/gpio_seqs.sv"
  
   `include "env_gpio/gpio_sequencer.sv"
   `include "env_gpio/gpio_driver.sv"
   `include "env_gpio/gpio_monitor.sv"
   `include "env_gpio/gpio_agent.sv"
  
   `include "env_gpio/axi_env.sv"
endpackage